--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:17:50 04/08/2018
-- Design Name:   
-- Module Name:   D:/Proyectos_Xilinx/Procesador1/test_UC.vhd
-- Project Name:  Procesador1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: UC
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY test_UC IS
END test_UC;
 
ARCHITECTURE behavior OF test_UC IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT UC
    PORT(
         entrada_OP : IN  std_logic_vector(1 downto 0);
         entrada_OP3 : IN  std_logic_vector(5 downto 0);
			SDR : out STD_LOGIC;
			WRENMEM: out STD_LOGIC;
			WRIN:out STD_LOGIC;
         salida_uc_op : OUT  std_logic_vector(5 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal entrada_OP : std_logic_vector(1 downto 0) := (others => '0');
   signal entrada_OP3 : std_logic_vector(5 downto 0) := (others => '0');

 	--Outputs
   signal salida_uc_op : std_logic_vector(5 downto 0);
	signal WRIN : STD_LOGIC;
	signal SDR :  STD_LOGIC;			
	signal WRENMEM: STD_LOGIC;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: UC PORT MAP (
          entrada_OP => entrada_OP,
          entrada_OP3 => entrada_OP3,
			 WRIN => WRIN,
			 SDR => SDR,
			 WRENMEM => WRENMEM,
          salida_uc_op => salida_uc_op
        );


 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		
		entrada_OP <= "10";
		entrada_OP3<="000100";
		
		
      wait for 100 ns;	

     -- wait for <clock>_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
